module iread_controller();
    


endmodule